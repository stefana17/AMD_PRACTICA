// Code your testbench here
// or browse Examples
module tb_siso;

  reg clkt;
  reg resett;
  reg sit;
  wire sot;
  
  //instantierea
  siso siso_inst(.clk(clkt),.reset(resett),.si(sit),.so(sot));

  //Generarea semnalului de ceas
  initial
    begin
		#0 clkt = 1'b0;
		forever #5 clkt = ~clkt;
	end

  initial 
    begin
    resett = 1; sit = 0;
    #10 resett = 0; // Dezactivarea semnalului de reset după 10 unități de timp
    #20 sit = 1; // Setarea si la 1 după 20 unități de timp
    #20 sit = 0; // Setarea si la 0 după alte 20 unități de timp
    end
  
  initial 
    begin
    #100 $finish; // Terminarea simulării după 100 unități de timp
    end
  
  initial
    begin
      $dumpfile("dump.vcd");
      $dumpvars(0, siso_inst);
    end

endmodule