module DataMemory(clk, we, address, writeData, readData);
  input clk, we;
  input address;
  output readData;
  reg [31:0] RAM [63:0];
  
  
endmodule
